-- mpultra_brd_decl
--
-- Defines constants for the whole device
--
-- Dave Newbold, June 2014

library IEEE;
use IEEE.STD_LOGIC_1164.all;

use work.emp_framework_decl;

-------------------------------------------------------------------------------
package mp7_top_decl is

  alias mgt_kind_t is work.emp_framework_decl.mgt_kind_t;
  alias chk_kind_t is work.emp_framework_decl.chk_kind_t;
  alias buf_kind_t is work.emp_framework_decl.buf_kind_t;
  alias fmt_kind_t is work.emp_framework_decl.fmt_kind_t;
  
end mp7_top_decl;
-------------------------------------------------------------------------------
